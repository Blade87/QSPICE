// Automatically generated .v file on Wed Feb 21 15:50:33 2024
//

module vlog ( in1, out1 ) ;
// You will probably want to flush out the nature of these port declarations:
   input real in1;
   output real out1;

   // Implement the module here
   assign out1 = in1 * in1 * in1;

endmodule
